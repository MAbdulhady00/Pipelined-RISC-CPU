module decode_exm_buffer ();
endmodule
